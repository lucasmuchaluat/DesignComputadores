library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 8;
          addrWidth: natural := 3
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
        -- Inicializa os endereços:
		  -- tmp -> OPCODE   Ra     Rb     Rc    IMEDIATO
				tmp(0):= b"01000000000011010000000000000001";
tmp(1):= b"01000000000001100000000000000000";
tmp(2):= b"01000000000010100000000000001001";
tmp(3):= b"01000000000010010000000000000101";
tmp(4):= b"01000000000001110000000000000010";
tmp(5):= b"01000000000011110000000000001000";
tmp(6):= b"01000000000010000000000000000011";
tmp(7):= b"10010000000000000000000000001000";
tmp(8):= b"01000000000011100000000000000000";
tmp(9):= b"01000000000001000000000000000000";
tmp(10):= b"01000000000001010000000000000000";
tmp(11):= b"01000000000000100000000000000000";
tmp(12):= b"01000000000000110000000000000000";
tmp(13):= b"01000000000000000000000000000000";
tmp(14):= b"01000000000000010000000000000000";
tmp(15):= b"10010000000000000000000000010000";
tmp(16):= b"01010100110100000000000000000000";
tmp(17):= b"10100000000000000000000000111001";
tmp(18):= b"10010000000000000000000000010011";
tmp(19):= b"00100001000000000000000000001110";
tmp(20):= b"00100000000000000000000000001111";
tmp(21):= b"00100010000000000000000000010001";
tmp(22):= b"00100011000000000000000000010000";
tmp(23):= b"00010000000010110000000000000010";
tmp(24):= b"01011101101100000000000000000000";
tmp(25):= b"10100000000000000000000000100010";
tmp(26):= b"10010000000000000000000000011011";
tmp(27):= b"00100101000000000000000000010010";
tmp(28):= b"00100100000000000000000000010011";
tmp(29):= b"10010000000000000000000000011110";
tmp(30):= b"00010000000010110000000000000011";
tmp(31):= b"01011101101100000000000000000000";
tmp(32):= b"10100000000000000000000000111110";
tmp(33):= b"10010000000000000000000001001101";
tmp(34):= b"00101110000000000000000000010100";
tmp(35):= b"01011110110100000000000000000000";
tmp(36):= b"10100000000000000000000000100110";
tmp(37):= b"10010000000000000000000000011011";
tmp(38):= b"01010100110100000000000000000000";
tmp(39):= b"10100000000000000000000000101001";
tmp(40):= b"10010000000000000000000000101101";
tmp(41):= b"00100110000000000000000000010011";
tmp(42):= b"10000101011110110000000000000000";
tmp(43):= b"00101011000000000000000000010010";
tmp(44):= b"10010000000000000000000000011110";
tmp(45):= b"01010101011000000000000000000000";
tmp(46):= b"10100000000000000000000000110101";
tmp(47):= b"01010101110100000000000000000000";
tmp(48):= b"10100000000000000000000000110101";
tmp(49):= b"00101101000000000000000000010011";
tmp(50):= b"10000101011110110000000000000000";
tmp(51):= b"00101011000000000000000000010010";
tmp(52):= b"10010000000000000000000000011110";
tmp(53):= b"00100110000000000000000000010011";
tmp(54):= b"01101111010110110000000000000000";
tmp(55):= b"00101011000000000000000000010010";
tmp(56):= b"10010000000000000000000000011110";
tmp(57):= b"01010101100000000000000000000000";
tmp(58):= b"10100000000000000000000000111100";
tmp(59):= b"10010000000000000000000000010011";
tmp(60):= b"01000000000011100000000000000001";
tmp(61):= b"10010000000000000000000000010011";
tmp(62):= b"00010000000010110000000000001000";
tmp(63):= b"01010110101100000000000000000000";
tmp(64):= b"10100000000000000000000001001001";
tmp(65):= b"00010000000010110000000000001001";
tmp(66):= b"01010110101100000000000000000000";
tmp(67):= b"10100000000000000000000001000101";
tmp(68):= b"10010000000000000000000000010011";
tmp(69):= b"00010000000010110000000000001001";
tmp(70):= b"01011101101100000000000000000000";
tmp(71):= b"10100000000000000000000001101001";
tmp(72):= b"10010000000000000000000001000101";
tmp(73):= b"00010000000010110000000000001000";
tmp(74):= b"01011101101100000000000000000000";
tmp(75):= b"10100000000000000000000001011101";
tmp(76):= b"10010000000000000000000001001001";
tmp(77):= b"00010000000011000000000000001100";
tmp(78):= b"01011101110000000000000000000000";
tmp(79):= b"10100000000000000000000001010001";
tmp(80):= b"10010000000000000000000000010000";
tmp(81):= b"00010000000011000000000000001101";
tmp(82):= b"01010001101000000000000000000000";
tmp(83):= b"10100000000000000000000001010111";
tmp(84):= b"01101101000110110000000000000000";
tmp(85):= b"00110000101100010000000000000000";
tmp(86):= b"10010000000000000000000000010000";
tmp(87):= b"00110000011000010000000000000000";
tmp(88):= b"01010000100100000000000000000000";
tmp(89):= b"10100000000000000000000001011101";
tmp(90):= b"01101101000010110000000000000000";
tmp(91):= b"00110000101100000000000000000000";
tmp(92):= b"10010000000000000000000000010000";
tmp(93):= b"00110000011000000000000000000000";
tmp(94):= b"01010011101000000000000000000000";
tmp(95):= b"10100000000000000000000001100011";
tmp(96):= b"01101101001110110000000000000000";
tmp(97):= b"00110000101100110000000000000000";
tmp(98):= b"10010000000000000000000000010000";
tmp(99):= b"00110000011000110000000000000000";
tmp(100):= b"01010010100100000000000000000000";
tmp(101):= b"10100000000000000000000001101001";
tmp(102):= b"01101101001010110000000000000000";
tmp(103):= b"00110000101100100000000000000000";
tmp(104):= b"10010000000000000000000000010000";
tmp(105):= b"00110000011000100000000000000000";
tmp(106):= b"01010101101000000000000000000000";
tmp(107):= b"10100000000000000000000001110001";
tmp(108):= b"01010101100000000000000000000000";
tmp(109):= b"10100000000000000000000001110101";
tmp(110):= b"01101101010110110000000000000000";
tmp(111):= b"00110000101101010000000000000000";
tmp(112):= b"10010000000000000000000000010000";
tmp(113):= b"00110000011001010000000000000000";
tmp(114):= b"01101101010010110000000000000000";
tmp(115):= b"00110000101101000000000000000000";
tmp(116):= b"10010000000000000000000000010000";
tmp(117):= b"01010100011100000000000000000000";
tmp(118):= b"10100000000000000000000000001000";
tmp(119):= b"10010000000000000000000001101110";
        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;